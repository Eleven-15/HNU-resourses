module psw(clk,cf_en,zf_en,cf,zf,c,z);
input clk,cf_en,zf_en,cf,zf;
output reg c,z;
always@(negedge clk)
begin
    if (cf_en) c<=cf;
    else c<=c;
    if (zf_en) z<=zf;
    else z<=z;
end
endmodule