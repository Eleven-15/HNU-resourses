library ieee;
use ieee.std_logic_1164.all;
entity xiuzheng is
port(
	cin:in std_logic_vector(3 downto 0);
	qa,qb,qc,qd,qe,qf,qg:in std_logic;
	qout:out std_logic_vector(6 downto 0));
end xiuzheng;

architecture exa of xiuzheng is
begin
	qout<=  "1110111"when cin ="1010"else
			"0011111"when cin ="1011"else
			"1001110"when cin ="1100"else
			"0111101"when cin ="1101"else
			"1001111"when cin ="1110"else
			"1000111"when cin ="1111"else
			qa&qb&qc&qd&qe&qf&qg;
end exa;
			